module pipelinedcpu(
    input wire clk,
    input wire start
);

