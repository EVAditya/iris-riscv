// module ifu( //Instruction fetch
//     input [6:0] opcode,  //Inst[6:0]
//     output  branch,
//     output  memRead,
//     output  memtoReg,
//     output  [1:0] ALUOp,
//     output  memWrite,
//     output  ALUSrc,
//     output  regWrite
// );

    
    
// endmodule